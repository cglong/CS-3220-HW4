library verilog;
use verilog.vl_types.all;
entity lg_highlevel is
end lg_highlevel;
